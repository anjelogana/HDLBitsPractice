//https://hdlbits.01xz.net/wiki/Step_one

module top_module( output one );

// Insert your code here
    assign one = 1'b1;

endmodule
