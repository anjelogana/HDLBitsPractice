https://hdlbits.01xz.net/wiki/Wire

module top_module( 
    input in, 
    output out);

    assign out = in;
    //Wires are Directional, assign in = out; is not a valid solution!
endmodule
